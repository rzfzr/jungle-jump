{"lastScore":0,"highScore":0,"totalScore":0,"tokens":1,"longestDistance":7,"longestStreak":3,"totalPowerups":0,"longestPowerUpStreak":0,"rounds":18}