{"lastScore":0,"highScore":0,"totalScore":0,"tokens":0,"longestDistance":14,"longestStreak":2,"totalPowerups":2,"longestPowerUpStreak":1,"rounds":7}