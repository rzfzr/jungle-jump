{"lastScore":0,"highScore":0,"totalScore":0,"tokens":0,"longestDistance":4,"longestStreak":1,"totalPowerups":0,"longestPowerUpStreak":0,"rounds":9}